module tb_draw();
    logic clock;
    logic rst_n;

endmodule